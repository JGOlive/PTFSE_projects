

module flsr(
        
    );

endmodule