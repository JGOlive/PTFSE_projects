`timescale 1ns / 1ps

module(
    input clk;
    input reset;
    input bist_start;
    input [1:0] in;
    output reg pass_nfail;
    output reg [1:0] out
    );



endmodule